module TOP();
endmodule
