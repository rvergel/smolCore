/*
	Author: Ricardo Vergel
	Description: COntrol module for smolCore datapath
	Date: April 22-2025
	
	****INSERT YOUR CHANGES BELOW****

*/

module smolControl(
	input logic [4:0] rd,
	input logic [31:0] imm,
	input logic [6:0] opcode,
	input logic [2:0] funct3,
	input logic funct7

	output [4:0] op_sel

);
endmodule
